module first (
    
);
initial begin
    $display("hello dip");
    $finish;
end
    
endmodule